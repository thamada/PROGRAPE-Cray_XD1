-------------------------------------------------------------------------------
-- Title      : RT Client
-- Project    : Hello World FPGA
-------------------------------------------------------------------------------
-- File       : $RCSfile: rt_client.vhd,v $
-- Author     : Cray Canada
-- Company    : Cray Canada Inc.
-- Created    : 2004-12-10
-- Last update: 2005-03-17
-------------------------------------------------------------------------------
-- Description: The RT Client block serves 'clients' of the RapidArray switch
-- fabric.  In other words, it handles the read and write requests generated by
-- other devices connected intended for the FPGA.  Currently, the only fabric
-- client is an Opteron processor.  In the case of the Opteron, this block
-- handles the requests generated when software on the Opteron makes calls
-- to the acceleration FPGA API.
-------------------------------------------------------------------------------
-- Copyright (c) 2004 Cray Canada Inc.
-------------------------------------------------------------------------------
-- Revisions  :
-- $Log: rt_client.vhd,v $
-- Revision 1.3  2005/03/17 19:54:20 
-- Changed the block_busy signal to two variables.
--
-- Revision 1.2  2005/01/25 22:48:08 
-- Changed some of the constant names.
--
-- Revision 1.1  2004/12/22 23:55:00 
-- Initial checkin.
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_misc.all;
use work.user_pkg.all;

entity rt_client is
  port (
    -- Global signals
    reset_n      : in  std_logic;
    user_clk     : in  std_logic;
    user_enable  : in  std_logic;
    rt_ready     : in  std_logic;
    -- RT Interface
    -- Fabric Request Interface
    freq_addr    : in  std_logic_vector(39 downto 3);  -- request address
    freq_size    : in  std_logic_vector(3 downto 0);   -- request size
    freq_mask    : in  std_logic_vector(7 downto 0);   -- request byte mask
    freq_rw_n    : in  std_logic;       -- request read/write 
    freq_ts      : in  std_logic;       -- request transfer start
    freq_valid   : in  std_logic;       -- request valid
    freq_data    : in  std_logic_vector(63 downto 0);  -- request write data
    freq_srctag  : in  std_logic_vector(4 downto 0);
    freq_enable  : out std_logic;       -- enable request interface
    -- User Response Interface
    uresp_full   : in  std_logic;       -- response buffer full
    uresp_ts     : out std_logic;       -- response transfer start
    uresp_size   : out std_logic_vector(3 downto 0);   -- response size
    uresp_data   : out std_logic_vector(63 downto 0);  -- response data
    uresp_srctag : out std_logic_vector(4 downto 0);   -- response source tag
    -- Block Interface
    rt_responses : in  t_rt_responses;
    rt_req       : out t_rt_req
    );

end entity rt_client;

architecture rtl of rt_client is

  -----------------------------------------------------------------------------
  -- Declare Types
  -----------------------------------------------------------------------------
  -- Declare a type for the request state machine.  This type defines the
  -- states of the state machine.
  type t_req_state is (idle, rd, rd_stall, wr, wr_stall);

  -- Declare an array of byte arrays so we can create 'pipelines' of registers.
  type t_data_array is array(t_rt_blocks) of t_byte_array(7 downto 0);

  -- Declare a record type to conveniently store fabric request information.
  type t_req_info is record
    ts     : std_logic;
    sel    : t_rt_sel;
    size   : std_logic_vector(3 downto 0);
    srctag : std_logic_vector(4 downto 0);
  end record t_req_info;

  -- Declare an array of these records so theat we can pipeline the request
  -- information. 
  type t_req_pipe is array(natural range <>) of t_req_info;

  -----------------------------------------------------------------------------
  -- Declare Constants
  -----------------------------------------------------------------------------

  -- Create an all zero info constant that can be used to reset any signals of
  -- type t_req_info.
  constant c_zero_info : t_req_info := (ts     => '0',
                                        sel    => (others => '0'),
                                        size   => (others => '0'),
                                        srctag => (others => '0'));

  constant c_req_delay  : natural := c_rt_block_max + 1;
  constant c_resp_delay : natural := c_rt_block_max + 1;

  -----------------------------------------------------------------------------
  -- Declare Components
  -----------------------------------------------------------------------------

  component delay is
    generic (
      no_cycles : natural); 
    port (
      clk      : in  std_logic;
      reset_n  : in  std_logic;
      data_in  : in  t_byte_array(7 downto 0);
      data_out : out t_byte_array(7 downto 0)); 
  end component delay;

  -----------------------------------------------------------------------------
  -- Declare Signals
  -----------------------------------------------------------------------------
  -- Fabric request signal registers.
  signal s_ts_r     : std_logic;
  signal s_rw_n_r   : std_logic;
  signal s_size_r   : std_logic_vector(3 downto 0);
  signal s_srctag_r : std_logic_vector(4 downto 0);
  signal s_ufull_r  : std_logic;
  signal s_addr_r   : std_logic_vector(39 downto 3);
  signal s_addr_r2  : std_logic_vector(39 downto 3);
  signal s_data_r   : t_byte_array(7 downto 0);
  signal s_data_r2  : t_byte_array(7 downto 0);
  signal s_mask_r   : std_logic_vector(7 downto 0);
  signal s_mask_r2  : std_logic_vector(7 downto 0);
  signal s_valid_r  : std_logic;
  signal s_valid_r2 : std_logic;
  
  -- Control signals
  signal s_req_state    : t_req_state;
  signal s_state_enable : std_logic;
  signal s_burst_count  : std_logic_vector(3 downto 0);
  signal s_freq_enable  : std_logic;

  -- Read Signals
  signal s_rd_req       : t_req_info;
  signal s_req_delay    : t_req_pipe(c_req_delay downto 0);
  signal s_data_delay   : t_data_array;
  signal s_uresp_data   : t_byte_array(7 downto 0);
  signal s_uresp_ts     : std_logic;
  signal s_uresp_size   : std_logic_vector(3 downto 0);
  signal s_uresp_srctag : std_logic_vector(4 downto 0);

  -- Block Interface Signals
  signal s_rt_req : t_rt_req;
  
begin  -- architecture rtl

  -----------------------------------------------------------------------------
  -- Fabric Request Input Registers
  -- This process latches the Fabric request signals for future use by the
  -- control logic and to drive the RAM outputs.
  -----------------------------------------------------------------------------
  freq_reg : process (user_clk, reset_n) is
  begin  -- process freq_reg
    if reset_n = '0' then               -- asynchronous reset (active low)
      s_valid_r      <= '0';
      s_addr_r       <= (others => '0');
      s_data_r       <= (others => (others => '0'));
      s_mask_r       <= (others => '0');
      s_rw_n_r       <= '0';
      s_valid_r2     <= '0';
      s_addr_r2      <= (others => '0');
      s_data_r2      <= (others => (others => '0'));
      s_mask_r2      <= (others => '0');
      s_size_r       <= (others => '0');
      s_ts_r         <= '0';
      s_srctag_r     <= (others => '0');
      s_state_enable <= '0';
    elsif user_clk'event and user_clk = '1' then  -- rising clock edge
      -- Fabric request input registers.
      -- These register latch all the fabric request signals to make
      -- it easier for the Xilinx tools to place the chip and still
      -- hit a high clock speed.  This is necessary since some of the signals
      -- have have high fan out.
      if (s_freq_enable = '1') then
        s_ts_r     <= freq_ts;
        s_size_r   <= freq_size;
        s_srctag_r <= freq_srctag;
        s_addr_r   <= freq_addr;
        s_rw_n_r   <= freq_rw_n;
        s_valid_r  <= freq_valid;
        s_valid_r2 <= s_valid_r;
        s_mask_r   <= freq_mask;
        s_mask_r2  <= s_mask_r;
        -- Assign each bit of the fabric request data bus to a byte_array type
        -- register so it can be manipulated more easily.
        for byte in 7 downto 0 loop
          s_data_r(byte) <= freq_data(byte*8+7 downto byte*8);
        end loop;  -- byte
        s_data_r2 <= s_data_r;
      end if;

      -- Load the address counter at the start of a request.  For the rest of
      -- the request, increment the bottom four bits for burst accesses.
      if (s_valid_r = '1' and s_ts_r = '1' and s_freq_enable = '1') then
        s_addr_r2 <= s_addr_r;
      elsif (s_req_state = rd or
             (s_req_state = wr and s_valid_r = '1')) then
        s_addr_r2(6 downto 3) <= s_addr_r2(6 downto 3) + 1;
      end if;

      -- Create an enable signal for the state machine.  Only enable the
      -- state machine when the user logic is ready (i.e. programmable clock
      -- is valid) and the RT Core is ready.
      s_state_enable <= user_enable and rt_ready;

    end if;
  end process freq_reg;

  -----------------------------------------------------------------------------
  -- Access Control.
  -- This process contains a state machine to generate the control signals
  -- necessary for read and write accesses.  It is controlled by the fabric
  -- request signals and a local burst transfer counter.
  -----------------------------------------------------------------------------
  access_control : process (user_clk, reset_n) is
    variable v_block_busy : std_logic;
    variable v_block_free : std_logic;
  begin  -- process access_control
    if reset_n = '0' then               -- asynchronous reset (active low)
      s_req_state   <= idle;
      s_freq_enable <= '0';
      s_burst_count <= (others => '0');
      s_ufull_r     <= '0';
    elsif user_clk'event and user_clk = '1' then        -- rising clock edge
      -- Set default values for the busy/free flags.
      v_block_busy := '0';
      v_block_free := '1';

      -- Create busy and free flags based on the target block's busy flag.
      for i in rt_responses'range loop
        if (s_addr_r(c_rt_block_match(i)'range) = c_rt_block_match(i)) then
          v_block_busy := rt_responses(i).busy;
        end if;
        if (s_addr_r2(c_rt_block_match(i)'range) = c_rt_block_match(i)) then
          v_block_free := not rt_responses(i).busy;
        end if;
      end loop;  -- i
      
      -- Register the user response full flag.  This makes the design a bit
      -- easier for the Xilinx tools to place.
      s_ufull_r <= uresp_full;
      
      -- Fabric request state machine.
      if (s_state_enable = '1') then
        case s_req_state is
          when idle =>
            if (s_ts_r = '1' and s_valid_r = '1') then  -- Valid start strobe.
              if (s_rw_n_r = '1') then  -- Start read.
                if (s_ufull_r = '0' or v_block_busy = '0') then
                  s_req_state <= rd;    -- Response buffer is free.
                else
                  s_req_state <= rd_stall;  -- Response is full so stall.
                end if;
                s_freq_enable <= '0';
              else                      -- Start write.
                if (v_block_busy = '1') then
                  s_req_state <= wr_stall;
                  s_freq_enable <= '0';
                else
                  s_req_state   <= wr;
                  s_freq_enable <= '1';
                end if;
              end if;
              s_burst_count <= s_size_r;
            else                        -- Sit on your butt.
              s_req_state   <= idle;
              s_burst_count <= (others => '0');
              s_freq_enable <= '1';
            end if;
          when rd =>
            case s_burst_count is
              when "0000" =>            -- Burst done. Go to idle.
                s_req_state   <= idle;
                s_freq_enable <= '1';
              when others =>            -- Continue burst read.
                s_req_state   <= rd;
                s_burst_count <= s_burst_count - 1;
                s_freq_enable <= '0';
            end case;
          when rd_stall =>              -- Wait on the response FIFO.
            if (s_ufull_r = '0' and v_block_free = '1') then
              s_req_state <= rd;
            else
              s_req_state <= rd_stall;
            end if;
            s_freq_enable <= '0';
          when wr =>
            case s_burst_count is
              when "0000" =>            -- Burst done.  Check for new request.
                if (s_ts_r = '1' and s_valid_r = '1') then
                  if (s_rw_n_r = '1') then  -- Start read.
                    if (s_ufull_r = '0') then
                      s_req_state <= rd;    -- Response buffer is free.
                    else
                      s_req_state <= rd_stall;  -- Response is full so stall.
                    end if;
                    s_freq_enable <= '0';
                  else                      -- Start write.
                    if (v_block_busy = '1') then
                      s_req_state <= wr_stall;
                      s_freq_enable <= '0';
                    else
                      s_req_state   <= wr;
                      s_freq_enable <= '1';
                    end if;
                  end if;
                  s_burst_count <= s_size_r;
                else                    -- Go to idle.
                  s_req_state   <= idle;
                  s_freq_enable <= '1';
                end if;
              when others =>            -- Continue burst write.
                s_req_state <= wr;
                if (s_valid_r = '1') then
                  s_burst_count <= s_burst_count - 1;
                end if;
                s_freq_enable <= '1';
            end case;
          when wr_stall =>              -- Wait on the block.
            if (v_block_free = '1') then
              s_req_state <= wr;
              s_freq_enable <= '1';
            else
              s_req_state <= wr_stall;
              s_freq_enable <= '0';
            end if;
          when others => null;
        end case;
      else -- Disabled.
        s_req_state   <= idle;
        s_freq_enable <= '0';
        s_burst_count <= (others => '0');
      end if;
    end if;
  end process access_control;

  -----------------------------------------------------------------------------
  -- RT Request
  -- Drive the rt_req bus that connects to other blocks in the design.
  -- For convenience, the fabric request information is re-packaged into a
  -- aggregate request signal that can be distibuted to the other blocks in the
  -- design.
  -----------------------------------------------------------------------------
  rt_request : process (user_clk, reset_n) is
  begin  -- process rt_request
    if reset_n = '0' then               -- asynchronous reset (active low)
      s_rt_req <= c_rt_req_zero;
    elsif user_clk'event and user_clk = '1' then  -- rising clock edge
      for i in t_rt_blocks loop
        if (s_addr_r2(c_rt_block_match(i)'range) = c_rt_block_match(i) and
            s_valid_r2 = '1' and s_req_state = wr) then
          s_rt_req.wr(i) <= '1';
        else
          s_rt_req.wr(i) <= '0';
        end if;
        if (s_addr_r2(c_rt_block_match(i)'range) = c_rt_block_match(i) and
            s_req_state = rd) then
          s_rt_req.rd(i) <= '1';
        else
          s_rt_req.rd(i) <= '0';
        end if;
      end loop;  -- i
      s_rt_req.addr  <= s_addr_r2(s_rt_req.addr'range);
      s_rt_req.mask  <= s_mask_r2;
      s_rt_req.wdata <= s_data_r2;
    end if;
  end process rt_request;

  -----------------------------------------------------------------------------
  -- Request Delay
  -- When requesting data from different blocks there is inevitably a latency
  -- between the time the request is issued and the time when the response data
  -- is available.  This process delays the request information long enough for
  -- the slowest device to respond.  The delayed information is then used to
  -- create the response.
  -----------------------------------------------------------------------------
  req_delay : process (user_clk, reset_n) is
  begin  -- process req_delay
    if (reset_n = '0') then
      s_rd_req    <= c_zero_info;
      s_req_delay <= (others => c_zero_info);
    elsif user_clk'event and user_clk = '1' then  -- rising clock edge
      -- Detect a read request and latch the request information.
      if (s_state_enable = '1' and s_valid_r = '1' and s_ts_r = '1' and
          s_freq_enable = '1') then
        s_rd_req.ts <= s_rw_n_r;
        for i in t_rt_blocks loop
          if (s_addr_r(c_rt_block_match(i)'range) = c_rt_block_match(i)) then
            s_rd_req.sel(i) <= '1';
          else
            s_rd_req.sel(i) <= '0';
          end if;
        end loop;  -- i
        s_rd_req.srctag <= s_srctag_r;
        s_rd_req.size   <= s_size_r;
      else
        s_rd_req.ts <= '0';
      end if;

      -- Put the request information into a pipeline do delay it.  The delayed
      -- information is used to generate a response at the appropriate time.
      s_req_delay(0).ts     <= s_rd_req.ts;
      s_req_delay(0).sel    <= s_rd_req.sel;
      s_req_delay(0).srctag <= s_rd_req.srctag;
      s_req_delay(0).size   <= s_rd_req.size;
      for stage in c_req_delay downto 1 loop
        s_req_delay(stage) <= s_req_delay(stage-1);
      end loop;  -- stage

    end if;
  end process req_delay;

  -----------------------------------------------------------------------------
  -- Response Delays
  -- Since responses from different blocks have different latency, variable
  -- delay registers are used to align the response data from different devices
  -- to the same point in time.  The delay block will generate a RAM based
  -- shift register to delay the data for the requested number of cycles.
  -----------------------------------------------------------------------------
  resp_delay_gen : for i in t_rt_blocks generate
    delay_inst : delay
      generic map (
        no_cycles => (c_resp_delay - c_rt_block_latency(i)))
      port map (
        clk      => user_clk,
        reset_n  => reset_n,
        data_in  => rt_responses(i).rdata,
        data_out => s_data_delay(i));
  end generate resp_delay_gen;
  
  -----------------------------------------------------------------------------
  -- RT User Response
  -- Create the signals required to drive the RT Core User Response bus.
  -- The user response signals are generated from the delayed request
  -- information.  The user response data is generated from the delayed
  -- data read in from the selected block.
  -----------------------------------------------------------------------------
  rt_resp : process (user_clk, reset_n) is
  begin  -- process rt_resp
    if reset_n = '0' then               -- asynchronous reset (active low)
      s_uresp_ts     <= '0';
      s_uresp_size   <= (others => '0');
      s_uresp_srctag <= (others => '0');
      s_uresp_data   <= (others => (others => '0'));
    elsif user_clk'event and user_clk = '1' then  -- rising clock edge
      -- Drive the response bus.
      s_uresp_ts     <= s_req_delay(c_req_delay).ts;
      s_uresp_size   <= s_req_delay(c_req_delay).size;
      s_uresp_srctag <= s_req_delay(c_req_delay).srctag;

      for i in t_rt_blocks loop
        if (s_req_delay(c_req_delay).sel(i) = '1') then
          s_uresp_data <= s_data_delay(i);
        end if;
      end loop;  -- i
    end if;
  end process rt_resp;


  -- Drive output ports with internal signals.
  freq_enable              <= s_freq_enable;

  uresp_data(7 downto 0)   <= s_uresp_data(0);
  uresp_data(15 downto 8)  <= s_uresp_data(1);
  uresp_data(23 downto 16) <= s_uresp_data(2);
  uresp_data(31 downto 24) <= s_uresp_data(3);
  uresp_data(39 downto 32) <= s_uresp_data(4);
  uresp_data(47 downto 40) <= s_uresp_data(5);
  uresp_data(55 downto 48) <= s_uresp_data(6);
  uresp_data(63 downto 56) <= s_uresp_data(7);

  uresp_ts                 <= s_uresp_ts;
  uresp_size               <= s_uresp_size;
  uresp_srctag             <= s_uresp_srctag;
  rt_req                   <= s_rt_req;

end architecture rtl;
